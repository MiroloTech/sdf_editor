module graph

// import os
// import x.json2 as json

/*
// TODO : Figure out compact structure
{
	"ui": {
		"panx": 20.0,
		"pany": 34.0,
		"dot_spacing": 50.0,
		"toast_lifetime": 4.0
	},
	"menu": {
		"math/simple": {
			"title": "Add",
			"pins": [
				"name": "A"
				
			]
		}
	}
}
*/


// Saves the graph in a specific structure as a .json file
pub fn (g Graph[T]) save(path string) ! {
	
}

pub fn (mut g Graph[T]) load(path string) ! {
	
}
